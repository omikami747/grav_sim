module interface (
                  );
endmodule
